module valida_rega(output [1:0]rega, output erro, input asp, input got, input [1:0] mef1, input limpeza);




endmodule
